LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Entit� du module de contr�le de la barri�re

ENTITY controle_barriere IS
  PORT (
    -- Signaux de contr�le
    clk   : IN  STD_LOGIC; -- Horloge (pour la logique s�quentielle)
    rst   : IN  STD_LOGIC; -- Reset asynchrone (pour initialiser)

    -- Entr�es (capteurs et commandes)
    trigger_open        : IN  STD_LOGIC; -- Ordre d'ouverture (vient du module principal)
    sensor_passage      : IN  STD_LOGIC; -- Capteur: la voiture est pass�e
    sensor_open_limit   : IN  STD_LOGIC; -- Capteur: la barri�re est en position haute
    sensor_closed_limit : IN  STD_LOGIC; -- Capteur: la barri�re est en position basse

    -- Sorties (commandes moteur)
    motor_open  : OUT STD_LOGIC; -- Commande au moteur: Ouvrir
    motor_close : OUT STD_LOGIC  -- Commande au moteur: Fermer
  );
END ENTITY controle_barriere;


-- Architecture 
-- Nous utilisons une machine � �tats (FSM)

ARCHITECTURE fsm OF controle_barriere IS

  -- 1. D�finition des �tats de notre FSM
  TYPE state_type IS (
    IDLE_CLOSED, -- La barri�re est ferm�e et attend
    OPENING,     -- La barri�re est en train de s'ouvrir
    IDLE_OPEN,   -- La barri�re est ouverte et attend le passage
    CLOSING      -- La barri�re est en train de se fermer
  );

  -- 2. Signal interne pour m�moriser l'�tat actuel et le prochain �tat
  SIGNAL state, next_state : state_type;

BEGIN

  -- PROCESS 1: Logique S�quentielle (Registre d'�tat)
  -- Ce process m�morise l'�tat actuel.
  -- Il est sensible au 'clk' et au 'rst', comme la bascule D (DFF)
  state_register_proc : PROCESS (clk, rst)
  BEGIN
    IF (rst = '1') THEN
      state <= IDLE_CLOSED; -- �tat initial de reset
    ELSIF (clk'EVENT AND clk = '1') THEN -- D�tection du front montant 
      state <= next_state; -- M�morisation du prochain �tat
    END IF;
  END PROCESS state_register_proc;


  -- PROCESS 2: Logique Combinatoire (Calcul du prochain �tat)
  -- Ce process calcule l'�tat suivant en fonction de l'�tat
  -- actuel et des entr�es (capteurs).
  next_state_logic_proc : PROCESS (state, trigger_open, sensor_passage, sensor_open_limit, sensor_closed_limit)
  BEGIN
    -- Par d�faut, on reste dans le m�me �tat
    next_state <= state; 

    CASE state IS
      -- �tat 1: Barri�re ferm�e
      WHEN IDLE_CLOSED =>
        IF (trigger_open = '1') THEN
          next_state <= OPENING; -- On passe � l'ouverture
        END IF;

      -- �tat 2: Barri�re en ouverture
      WHEN OPENING =>
        IF (sensor_open_limit = '1') THEN
          next_state <= IDLE_OPEN; -- On est arriv� en haut
        END IF;

      -- �tat 3: Barri�re ouverte
      WHEN IDLE_OPEN =>
        IF (sensor_passage = '1') THEN
          next_state <= CLOSING; -- La voiture est pass�e, on ferme
        END IF;

      -- �tat 4: Barri�re en fermeture
      WHEN CLOSING =>
        IF (sensor_closed_limit = '1') THEN
          next_state <= IDLE_CLOSED; -- On est arriv� en bas, retour � l'�tat initial
        END IF;

      -- Cas par d�faut (s�curit�)
      WHEN OTHERS =>
        next_state <= IDLE_CLOSED;

    END CASE;
  END PROCESS next_state_logic_proc;


  -- PROCESS 3: Logique Combinatoire (Logique de sortie)
  -- Ce process d�termine les sorties (commandes moteur)
  -- en fonction de l'�tat actuel.
  output_logic_proc : PROCESS (state)
  BEGIN
    -- Valeurs par d�faut pour �viter les "latches"
    motor_open  <= '0';
    motor_close <= '0';

    CASE state IS
      WHEN IDLE_CLOSED =>
        motor_open  <= '0';
        motor_close <= '0';
      
      WHEN OPENING =>
        motor_open  <= '1'; -- On active le moteur pour ouvrir
        motor_close <= '0';
      
      WHEN IDLE_OPEN =>
        motor_open  <= '0';
        motor_close <= '0';
      
      WHEN CLOSING =>
        motor_open  <= '0';
        motor_close <= '1'; -- On active le moteur pour fermer
      
      WHEN OTHERS =>
        motor_open  <= '0';
        motor_close <= '0';
        
    END CASE;
  END PROCESS output_logic_proc;

END ARCHITECTURE fsm;
