LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- L'entit� du testbench
ENTITY tb_controle_barriere IS
END ENTITY tb_controle_barriere;


ARCHITECTURE test OF tb_controle_barriere IS

  -- 1. D�clarer le composant � tester (votre module)
  COMPONENT controle_barriere
    PORT (
      clk                   : IN  STD_LOGIC;
      rst                   : IN  STD_LOGIC;
      trigger_open        : IN  STD_LOGIC;
      sensor_passage      : IN  STD_LOGIC;
      sensor_open_limit   : IN  STD_LOGIC;
      sensor_closed_limit : IN  STD_LOGIC;
      motor_open          : OUT STD_LOGIC;
      motor_close         : OUT STD_LOGIC
    );
  END COMPONENT;

  -- 2. Cr�er les signaux pour se connecter au composant
  -- Signaux d'entr�e (stimuli)
  SIGNAL s_clk                 : STD_LOGIC := '0';
  SIGNAL s_rst                 : STD_LOGIC;
  SIGNAL s_trigger_open        : STD_LOGIC := '0';
  SIGNAL s_sensor_passage      : STD_LOGIC := '0';
  SIGNAL s_sensor_open_limit   : STD_LOGIC := '0';
  SIGNAL s_sensor_closed_limit : STD_LOGIC := '0';

  -- Signaux de sortie (observation)
  SIGNAL s_motor_open  : STD_LOGIC;
  SIGNAL s_motor_close : STD_LOGIC;

  -- P�riode d'horloge
  CONSTANT CLK_PERIOD : TIME := 10 ns; -- Horloge de 100 MHz

BEGIN

  -- 3. Instancier le DUT (Device Under Test)
  -- On connecte les signaux du testbench aux ports du module
  DUT : controle_barriere
    PORT MAP (
      clk                   => s_clk,
      rst                   => s_rst,
      trigger_open        => s_trigger_open,
      sensor_passage      => s_sensor_passage,
      sensor_open_limit   => s_sensor_open_limit,
      sensor_closed_limit => s_sensor_closed_limit,
      motor_open          => s_motor_open,
      motor_close         => s_motor_close
    );

  -- 4. G�n�rateur d'horloge 
  clk_gen_proc : PROCESS
  BEGIN
    s_clk <= '0';
    WAIT FOR CLK_PERIOD / 2;
    s_clk <= '1';
    WAIT FOR CLK_PERIOD / 2;
  END PROCESS clk_gen_proc;


  -- 5. Processus de simulation (sc�nario de test)
  stimulus_proc : PROCESS
  BEGIN
    -- == PHASE 1: RESET ==
    s_rst <= '1'; -- Appliquer le reset
    WAIT FOR 20 ns;
    s_rst <= '0'; -- Rel�cher le reset
    WAIT FOR 10 ns;
    -- � ce stade, la FSM doit �tre dans l'�tat IDLE_CLOSED
    -- et les moteurs doivent �tre � '0'.

    -- == PHASE 2: SC�NARIO D'OUVERTURE ==
    s_trigger_open <= '1'; -- Le module principal demande l'ouverture
    WAIT FOR CLK_PERIOD;
    s_trigger_open <= '0'; -- L'ordre est une impulsion
    
    -- La FSM doit passer � OPENING. s_motor_open doit passer � '1'.
    WAIT FOR 50 ns; -- Simule le temps que prend la barri�re pour s'ouvrir

    -- Le capteur de limite haute est atteint
    s_sensor_open_limit <= '1';
    WAIT FOR CLK_PERIOD;
    s_sensor_open_limit <= '0';
    
    -- La FSM doit passer � IDLE_OPEN. Les moteurs doivent s'arr�ter.
    WAIT FOR 100 ns; -- Simule la voiture qui passe sous la barri�re

    -- == PHASE 3: SC�NARIO DE FERMETURE ==
    -- La voiture a activ� le capteur de passage
    s_sensor_passage <= '1';
    WAIT FOR CLK_PERIOD;
    s_sensor_passage <= '0';

    -- La FSM doit passer � CLOSING. s_motor_close doit passer � '1'.
    WAIT FOR 50 ns; -- Simule le temps que prend la barri�re pour se fermer

    -- Le capteur de limite basse est atteint
    s_sensor_closed_limit <= '1';
    WAIT FOR CLK_PERIOD;
    s_sensor_closed_limit <= '0';
    
    -- La FSM doit revenir � IDLE_CLOSED. Les moteurs doivent s'arr�ter.

    -- == FIN DE LA SIMULATION ==
    WAIT; 
  END PROCESS stimulus_proc;

END ARCHITECTURE test;
